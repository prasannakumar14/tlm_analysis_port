package pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;

  `include "xtn.sv"
  `include "producer.sv"
  `include "consumer.sv"
  `include "env.sv"
  `include "test.sv"
endpackage
